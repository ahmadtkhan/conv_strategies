// dsp.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module dsp (
		input  wire [1:0]  aclr,    //    aclr.aclr
		input  wire [17:0] ax,      //      ax.ax
		input  wire [17:0] ay,      //      ay.ay
		input  wire [17:0] bx,      //      bx.bx
		input  wire [17:0] by,      //      by.by
		input  wire [2:0]  clk,     //     clk.clk
		input  wire [2:0]  ena,     //     ena.ena
		output wire [36:0] resulta, // resulta.resulta
		output wire [36:0] resultb  // resultb.resultb
	);

	dsp_altera_a10_native_fixed_point_dsp_201_ffpppjq a10_native_fixed_point_dsp_0 (
		.ay      (ay),      //      ay.ay
		.by      (by),      //      by.by
		.ax      (ax),      //      ax.ax
		.bx      (bx),      //      bx.bx
		.resulta (resulta), // resulta.resulta
		.resultb (resultb), // resultb.resultb
		.clk     (clk),     //     clk.clk
		.ena     (ena),     //     ena.ena
		.aclr    (aclr)     //    aclr.aclr
	);

endmodule
